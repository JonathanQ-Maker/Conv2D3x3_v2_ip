`ifndef DEFINITIONS
`define DEFINITIONS

`define WORD_WIDTH 8
`define MAX_DEPTH 10

`endif