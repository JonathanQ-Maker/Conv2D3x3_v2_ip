`ifndef DEFINITIONS
`define DEFINITIONS

`define WIDTH 8
`define MAX_DEPTH 3

`endif