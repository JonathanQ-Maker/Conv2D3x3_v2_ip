`ifndef DEFINITIONS
`define DEFINITIONS

`define WORD_WIDTH 8
`define MAX_IMG_WIDTH 6
`define MAX_IMG_HEIGHT 6
`define MAX_TRANSFERS 3

`endif