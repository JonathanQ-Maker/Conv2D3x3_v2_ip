`ifndef DEFINITIONS
`define DEFINITIONS

`define TRANSFER_WIDTH 8
`define WORD_WIDTH 8

`define MAX_IMG_WIDTH 128
`define MAX_IMG_HEIGHT 128
`define MAX_TRANSFERS 3

`define MAX_LINE_DEPTH 8192
`define MAX_KERNEL_DEPTH 8
`define ADDR_WIDTH 32

`endif