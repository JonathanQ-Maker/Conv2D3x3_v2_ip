`ifndef DEFINITIONS
`define DEFINITIONS

`define WORD_WIDTH 8
`define NUM_TERMS 9

`endif