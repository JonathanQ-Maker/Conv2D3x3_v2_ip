`ifndef DEFINITIONS
`define DEFINITIONS

`define TRANSFER_WIDTH 8
`define WORD_WIDTH 8
`define MAX_FILTERS 6
`define MAX_TRANSFERS 3


`endif